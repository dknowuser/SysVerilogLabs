// qlab5_sys_tb.v

// Generated using ACDS version 12.1sp1 243 at 2020.03.08.17:33:30

`timescale 1 ps / 1 ps
module qlab5_sys_tb (
	);

	wire    qlab5_sys_inst_clk_0_clk_in_bfm_clk_clk;           // qlab5_sys_inst_clk_0_clk_in_bfm:clk -> [qlab5_sys_inst:clk_0, qlab5_sys_inst_clk_0_clk_in_reset_bfm:clk]
	wire    qlab5_sys_inst_clk_0_clk_in_reset_bfm_reset_reset; // qlab5_sys_inst_clk_0_clk_in_reset_bfm:reset -> qlab5_sys_inst:reset_n

	qlab5_sys qlab5_sys_inst (
		.clk_0                   (qlab5_sys_inst_clk_0_clk_in_bfm_clk_clk),           //              clk_0_clk_in.clk
		.reset_n                 (qlab5_sys_inst_clk_0_clk_in_reset_bfm_reset_reset), //        clk_0_clk_in_reset.reset_n
		.out_port_from_the_pio_0 ()                                                   // pio_0_external_connection.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) qlab5_sys_inst_clk_0_clk_in_bfm (
		.clk (qlab5_sys_inst_clk_0_clk_in_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) qlab5_sys_inst_clk_0_clk_in_reset_bfm (
		.reset (qlab5_sys_inst_clk_0_clk_in_reset_bfm_reset_reset), // reset.reset_n
		.clk   (qlab5_sys_inst_clk_0_clk_in_bfm_clk_clk)            //   clk.clk
	);

endmodule
