library verilog;
use verilog.vl_types.all;
entity \bus\ is
end \bus\;
