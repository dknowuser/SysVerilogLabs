library verilog;
use verilog.vl_types.all;
entity test_st_m is
end test_st_m;
