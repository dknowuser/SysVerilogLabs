library verilog;
use verilog.vl_types.all;
entity Test_sv is
end Test_sv;
