// flab5_tb.v

// Generated using ACDS version 12.1sp1 243 at 2020.03.08.21:25:28

`timescale 1 ps / 1 ps
module flab5_tb (
	);

	wire        flab5_inst_clk_bfm_clk_clk;       // flab5_inst_clk_bfm:clk -> [flab5_inst:clk_clk, flab5_inst_reset_bfm:clk]
	wire        flab5_inst_reset_bfm_reset_reset; // flab5_inst_reset_bfm:reset -> flab5_inst:reset_reset_n
	wire  [7:0] flab5_inst_out_data_export;       // flab5_inst:out_data_export -> flab5_inst_out_data_bfm:sig_export

	flab5 flab5_inst (
		.clk_clk         (flab5_inst_clk_bfm_clk_clk),       //      clk.clk
		.reset_reset_n   (flab5_inst_reset_bfm_reset_reset), //    reset.reset_n
		.out_data_export (flab5_inst_out_data_export)        // out_data.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) flab5_inst_clk_bfm (
		.clk (flab5_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) flab5_inst_reset_bfm (
		.reset (flab5_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (flab5_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm flab5_inst_out_data_bfm (
		.sig_export (flab5_inst_out_data_export)  // conduit.export
	);

endmodule
