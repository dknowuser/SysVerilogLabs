library verilog;
use verilog.vl_types.all;
entity altera_mult_add_rtl is
    generic(
        extra_latency   : integer := 0;
        dedicated_multiplier_circuitry: string  := "AUTO";
        dsp_block_balancing: string  := "AUTO";
        selected_device_family: string  := "Stratix V";
        lpm_type        : string  := "altmult_add";
        lpm_hint        : string  := "UNUSED";
        width_a         : integer := 1;
        input_register_a0: string  := "UNREGISTERED";
        input_aclr_a0   : string  := "NONE";
        input_source_a0 : string  := "DATAA";
        input_register_a1: string  := "UNREGISTERED";
        input_aclr_a1   : string  := "NONE";
        input_source_a1 : string  := "DATAA";
        input_register_a2: string  := "UNREGISTERED";
        input_aclr_a2   : string  := "NONE";
        input_source_a2 : string  := "DATAA";
        input_register_a3: string  := "UNREGISTERED";
        input_aclr_a3   : string  := "NONE";
        input_source_a3 : string  := "DATAA";
        width_b         : integer := 1;
        input_register_b0: string  := "UNREGISTERED";
        input_aclr_b0   : string  := "NONE";
        input_source_b0 : string  := "DATAB";
        input_register_b1: string  := "UNREGISTERED";
        input_aclr_b1   : string  := "NONE";
        input_source_b1 : string  := "DATAB";
        input_register_b2: string  := "UNREGISTERED";
        input_aclr_b2   : string  := "NONE";
        input_source_b2 : string  := "DATAB";
        input_register_b3: string  := "UNREGISTERED";
        input_aclr_b3   : string  := "NONE";
        input_source_b3 : string  := "DATAB";
        width_c         : integer := 1;
        input_register_c0: string  := "UNREGISTERED";
        input_aclr_c0   : string  := "NONE";
        input_register_c1: string  := "UNREGISTERED";
        input_aclr_c1   : string  := "NONE";
        input_register_c2: string  := "UNREGISTERED";
        input_aclr_c2   : string  := "NONE";
        input_register_c3: string  := "UNREGISTERED";
        input_aclr_c3   : string  := "NONE";
        width_result    : integer := 34;
        output_register : string  := "UNREGISTERED";
        output_aclr     : string  := "NONE";
        port_signa      : string  := "PORT_UNUSED";
        representation_a: string  := "UNSIGNED";
        signed_register_a: string  := "UNREGISTERED";
        signed_aclr_a   : string  := "NONE";
        signed_pipeline_register_a: string  := "UNREGISTERED";
        signed_pipeline_aclr_a: string  := "NONE";
        port_signb      : string  := "PORT_UNUSED";
        representation_b: string  := "UNSIGNED";
        signed_register_b: string  := "UNREGISTERED";
        signed_aclr_b   : string  := "NONE";
        signed_pipeline_register_b: string  := "UNREGISTERED";
        signed_pipeline_aclr_b: string  := "NONE";
        number_of_multipliers: integer := 1;
        multiplier1_direction: string  := "NONE";
        multiplier3_direction: string  := "NONE";
        multiplier_register0: string  := "UNREGISTERED";
        multiplier_aclr0: string  := "NONE";
        multiplier_register1: string  := "UNREGISTERED";
        multiplier_aclr1: string  := "NONE";
        multiplier_register2: string  := "UNREGISTERED";
        multiplier_aclr2: string  := "NONE";
        multiplier_register3: string  := "UNREGISTERED";
        multiplier_aclr3: string  := "NONE";
        port_addnsub1   : string  := "PORT_UNUSED";
        addnsub_multiplier_register1: string  := "UNREGISTERED";
        addnsub_multiplier_aclr1: string  := "NONE";
        addnsub_multiplier_pipeline_register1: string  := "UNREGISTERED";
        addnsub_multiplier_pipeline_aclr1: string  := "NONE";
        port_addnsub3   : string  := "PORT_UNUSED";
        addnsub_multiplier_register3: string  := "UNREGISTERED";
        addnsub_multiplier_aclr3: string  := "NONE";
        addnsub_multiplier_pipeline_register3: string  := "UNREGISTERED";
        addnsub_multiplier_pipeline_aclr3: string  := "NONE";
        adder1_rounding : string  := "NO";
        addnsub1_round_register: string  := "UNREGISTERED";
        addnsub1_round_aclr: string  := "NONE";
        addnsub1_round_pipeline_register: string  := "UNREGISTERED";
        addnsub1_round_pipeline_aclr: string  := "NONE";
        adder3_rounding : string  := "NO";
        addnsub3_round_register: string  := "UNREGISTERED";
        addnsub3_round_aclr: string  := "NONE";
        addnsub3_round_pipeline_register: string  := "UNREGISTERED";
        addnsub3_round_pipeline_aclr: string  := "NONE";
        multiplier01_rounding: string  := "NO";
        mult01_round_register: string  := "UNREGISTERED";
        mult01_round_aclr: string  := "NONE";
        multiplier23_rounding: string  := "NO";
        mult23_round_register: string  := "UNREGISTERED";
        mult23_round_aclr: string  := "NONE";
        width_msb       : integer := 17;
        output_rounding : string  := "NO";
        output_round_type: string  := "NEAREST_INTEGER";
        output_round_register: string  := "UNREGISTERED";
        output_round_aclr: string  := "NONE";
        output_round_pipeline_register: string  := "UNREGISTERED";
        output_round_pipeline_aclr: string  := "NONE";
        chainout_rounding: string  := "NO";
        chainout_round_register: string  := "UNREGISTERED";
        chainout_round_aclr: string  := "NONE";
        chainout_round_pipeline_register: string  := "UNREGISTERED";
        chainout_round_pipeline_aclr: string  := "NONE";
        chainout_round_output_register: string  := "UNREGISTERED";
        chainout_round_output_aclr: string  := "NONE";
        multiplier01_saturation: string  := "NO";
        mult01_saturation_register: string  := "UNREGISTERED";
        mult01_saturation_aclr: string  := "NONE";
        multiplier23_saturation: string  := "NO";
        mult23_saturation_register: string  := "UNREGISTERED";
        mult23_saturation_aclr: string  := "NONE";
        port_mult0_is_saturated: string  := "NONE";
        port_mult1_is_saturated: string  := "NONE";
        port_mult2_is_saturated: string  := "NONE";
        port_mult3_is_saturated: string  := "NONE";
        width_saturate_sign: integer := 1;
        output_saturation: string  := "NO";
        port_output_is_overflow: string  := "PORT_UNUSED";
        output_saturate_type: string  := "ASYMMETRIC";
        output_saturate_register: string  := "UNREGISTERED";
        output_saturate_aclr: string  := "NONE";
        output_saturate_pipeline_register: string  := "UNREGISTERED";
        output_saturate_pipeline_aclr: string  := "NONE";
        chainout_saturation: string  := "NO";
        port_chainout_sat_is_overflow: string  := "PORT_UNUSED";
        chainout_saturate_register: string  := "UNREGISTERED";
        chainout_saturate_aclr: string  := "NONE";
        chainout_saturate_pipeline_register: string  := "UNREGISTERED";
        chainout_saturate_pipeline_aclr: string  := "NONE";
        chainout_saturate_output_register: string  := "UNREGISTERED";
        chainout_saturate_output_aclr: string  := "NONE";
        scanouta_register: string  := "UNREGISTERED";
        scanouta_aclr   : string  := "NONE";
        width_chainin   : integer := 1;
        chainout_adder  : string  := "NO";
        chainout_register: string  := "UNREGISTERED";
        chainout_aclr   : string  := "NONE";
        zero_chainout_output_register: string  := "UNREGISTERED";
        zero_chainout_output_aclr: string  := "NONE";
        shift_mode      : string  := "NO";
        rotate_register : string  := "UNREGISTERED";
        rotate_aclr     : string  := "NONE";
        rotate_pipeline_register: string  := "UNREGISTERED";
        rotate_pipeline_aclr: string  := "NONE";
        rotate_output_register: string  := "UNREGISTERED";
        rotate_output_aclr: string  := "NONE";
        shift_right_register: string  := "UNREGISTERED";
        shift_right_aclr: string  := "NONE";
        shift_right_pipeline_register: string  := "UNREGISTERED";
        shift_right_pipeline_aclr: string  := "NONE";
        shift_right_output_register: string  := "UNREGISTERED";
        shift_right_output_aclr: string  := "NONE";
        zero_loopback_register: string  := "UNREGISTERED";
        zero_loopback_aclr: string  := "NONE";
        zero_loopback_pipeline_register: string  := "UNREGISTERED";
        zero_loopback_pipeline_aclr: string  := "NONE";
        zero_loopback_output_register: string  := "UNREGISTERED";
        zero_loopback_output_aclr: string  := "NONE";
        accumulator     : string  := "NO";
        accum_direction : string  := "ADD";
        loadconst_value : integer := 0;
        use_sload_accum_port: string  := "NO";
        accum_sload_register: string  := "UNREGISTERED";
        accum_sload_aclr: string  := "NONE";
        accum_sload_pipeline_register: string  := "UNREGISTERED";
        accum_sload_pipeline_aclr: string  := "NONE";
        loadconst_control_register: string  := "UNREGISTERED";
        loadconst_control_aclr: string  := "NONE";
        double_accum    : string  := "NO";
        systolic_delay1 : string  := "UNREGISTERED";
        systolic_delay3 : string  := "UNREGISTERED";
        systolic_aclr1  : string  := "NONE";
        systolic_aclr3  : string  := "NONE";
        preadder_mode   : string  := "SIMPLE";
        preadder_direction_0: string  := "ADD";
        preadder_direction_1: string  := "ADD";
        preadder_direction_2: string  := "ADD";
        preadder_direction_3: string  := "ADD";
        width_coef      : integer := 1;
        coefsel0_register: string  := "UNREGISTERED";
        coefsel0_aclr   : string  := "NONE";
        coefsel1_register: string  := "UNREGISTERED";
        coefsel1_aclr   : string  := "NONE";
        coefsel2_register: string  := "UNREGISTERED";
        coefsel2_aclr   : string  := "NONE";
        coefsel3_register: string  := "UNREGISTERED";
        coefsel3_aclr   : string  := "NONE";
        coef0_0         : integer := 0;
        coef0_1         : integer := 0;
        coef0_2         : integer := 0;
        coef0_3         : integer := 0;
        coef0_4         : integer := 0;
        coef0_5         : integer := 0;
        coef0_6         : integer := 0;
        coef0_7         : integer := 0;
        coef1_0         : integer := 0;
        coef1_1         : integer := 0;
        coef1_2         : integer := 0;
        coef1_3         : integer := 0;
        coef1_4         : integer := 0;
        coef1_5         : integer := 0;
        coef1_6         : integer := 0;
        coef1_7         : integer := 0;
        coef2_0         : integer := 0;
        coef2_1         : integer := 0;
        coef2_2         : integer := 0;
        coef2_3         : integer := 0;
        coef2_4         : integer := 0;
        coef2_5         : integer := 0;
        coef2_6         : integer := 0;
        coef2_7         : integer := 0;
        coef3_0         : integer := 0;
        coef3_1         : integer := 0;
        coef3_2         : integer := 0;
        coef3_3         : integer := 0;
        coef3_4         : integer := 0;
        coef3_5         : integer := 0;
        coef3_6         : integer := 0;
        coef3_7         : integer := 0;
        width_clock_all_wire_msb: integer := 3;
        width_aclr_all_wire_msb: integer := 3;
        width_ena_all_wire_msb: integer := 3
    );
    port(
        dataa           : in     vl_logic_vector;
        datab           : in     vl_logic_vector;
        datac           : in     vl_logic_vector;
        scanina         : in     vl_logic_vector;
        scaninb         : in     vl_logic_vector;
        sourcea         : in     vl_logic_vector;
        sourceb         : in     vl_logic_vector;
        clock3          : in     vl_logic;
        clock2          : in     vl_logic;
        clock1          : in     vl_logic;
        clock0          : in     vl_logic;
        aclr3           : in     vl_logic;
        aclr2           : in     vl_logic;
        aclr1           : in     vl_logic;
        aclr0           : in     vl_logic;
        ena3            : in     vl_logic;
        ena2            : in     vl_logic;
        ena1            : in     vl_logic;
        ena0            : in     vl_logic;
        signa           : in     vl_logic;
        signb           : in     vl_logic;
        addnsub1        : in     vl_logic;
        addnsub3        : in     vl_logic;
        result          : out    vl_logic_vector;
        scanouta        : out    vl_logic_vector;
        scanoutb        : out    vl_logic_vector;
        mult01_round    : in     vl_logic;
        mult23_round    : in     vl_logic;
        mult01_saturation: in     vl_logic;
        mult23_saturation: in     vl_logic;
        addnsub1_round  : in     vl_logic;
        addnsub3_round  : in     vl_logic;
        mult0_is_saturated: out    vl_logic;
        mult1_is_saturated: out    vl_logic;
        mult2_is_saturated: out    vl_logic;
        mult3_is_saturated: out    vl_logic;
        output_round    : in     vl_logic;
        chainout_round  : in     vl_logic;
        output_saturate : in     vl_logic;
        chainout_saturate: in     vl_logic;
        overflow        : out    vl_logic;
        chainout_sat_overflow: out    vl_logic;
        chainin         : in     vl_logic_vector;
        zero_chainout   : in     vl_logic;
        rotate          : in     vl_logic;
        shift_right     : in     vl_logic;
        zero_loopback   : in     vl_logic;
        accum_sload     : in     vl_logic;
        sload_accum     : in     vl_logic;
        coefsel0        : in     vl_logic_vector(2 downto 0);
        coefsel1        : in     vl_logic_vector(2 downto 0);
        coefsel2        : in     vl_logic_vector(2 downto 0);
        coefsel3        : in     vl_logic_vector(2 downto 0)
    );
end altera_mult_add_rtl;
