/*module flab5(input wire clk, input wire reset_n,
	output wire data_out);

flab5_sys flab5_cpu(.clk_0(clk), .reset_n(reset_n),
	.out_port_from_the_pio_0(data_out));

endmodule*/